/***********************************************
Module Name:   square_read_create_test
Feature:       Testbench for square_read_create
               An example for the book
Coder:         Garfield
Organization:  XXXX Group, Department of Architecture
------------------------------------------------------
Variables:
         clk: clock for processing
         reset: reset flag
----------------------------------------------------
History:
03-01-2016: First Version by Garfield
***********************************************/
`timescale 10 ns/100 ps
//Simulation time assignment

//Insert the modules

module square_read_create_test;
//defination for Variables
reg clk;
reg reset;

reg[5:0] counter;
wire[11:0] square_file, square;

//Connection to the modules
square_read_create C1( .CLK(clk), .RST(reset),
 	  .square(square_file) );

begin

assign square = counter * counter;
 
//Clock generation
    initial
    begin
      clk = 0;
      //Reset
      forever  
      begin
           #10 clk = !clk;
           //Reverse the clock in each 10ns
      end
    end

//Reset operation
    initial  
    begin
      reset = 0;
      //Reset enable
      #14  reset = 1;
     //Counter starts
    end
end

always @(posedge clk or negedge reset)
//Counter
begin
    if ( !reset)
    begin
        counter <= 6'h00;
        //Reset
    end
    else
    begin
        counter <= counter + 6'h01;
        //Increase
    end
end
endmodule